module HexHELO(Hex, C);
	input [2:0] C;
	output [0:6] Hex;
	
	assign Seg
	
endmodule	